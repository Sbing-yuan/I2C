module DLY_chain(
    IN,
    D80,
);

input   IN;
output  D80;

lcell  U0(.in(IN)    , .out(SD1));
lcell  U1(.in(SD1)   , .out(SD2));
lcell  U2(.in(SD2)   , .out(SD3));
lcell  U3(.in(SD3)   , .out(SD4));
lcell  U4(.in(SD4)   , .out(SD5));
lcell  U5(.in(SD5)   , .out(SD6));
lcell  U6(.in(SD6)   , .out(SD7));
lcell  U7(.in(SD7)   , .out(SD8));
lcell  U8(.in(SD8)   , .out(SD9));
lcell  U9(.in(SD9)   , .out(SD10));
lcell U10(.in(SD10)  , .out(SD11));
lcell U11(.in(SD11)  , .out(SD12));
lcell U12(.in(SD12)  , .out(SD13));
lcell U13(.in(SD13)  , .out(SD14));
lcell U14(.in(SD14)  , .out(SD15));
lcell U15(.in(SD15)  , .out(SD16));
lcell U16(.in(SD16)  , .out(SD17));
lcell U17(.in(SD17)  , .out(SD18));
lcell U18(.in(SD18)  , .out(SD19));
lcell U19(.in(SD19)  , .out(SD20));
lcell U20(.in(SD20)  , .out(SD21));
lcell U21(.in(SD21)  , .out(SD22));
lcell U22(.in(SD22)  , .out(SD23));
lcell U23(.in(SD23)  , .out(SD24));
lcell U24(.in(SD24)  , .out(SD25));
lcell U25(.in(SD25)  , .out(SD26));
lcell U26(.in(SD26)  , .out(SD27));
lcell U27(.in(SD27)  , .out(SD28));
lcell U28(.in(SD28)  , .out(SD29));
lcell U29(.in(SD29)  , .out(SD30));
lcell U30(.in(SD30)  , .out(SD31));
lcell U31(.in(SD31)  , .out(SD32));
lcell U32(.in(SD32)  , .out(SD33));
lcell U33(.in(SD33)  , .out(SD34));
lcell U34(.in(SD34)  , .out(SD35));
lcell U35(.in(SD35)  , .out(SD36));
lcell U36(.in(SD36)  , .out(SD37));
lcell U37(.in(SD37)  , .out(SD38));
lcell U38(.in(SD38)  , .out(SD39));
lcell U39(.in(SD39)  , .out(SD40));
lcell U40(.in(SD40)  , .out(SD41));
lcell U41(.in(SD41)  , .out(SD42));
lcell U42(.in(SD42)  , .out(SD43));
lcell U43(.in(SD43)  , .out(SD44));
lcell U44(.in(SD44)  , .out(SD45));
lcell U45(.in(SD45)  , .out(SD46));
lcell U46(.in(SD46)  , .out(SD47));
lcell U47(.in(SD47)  , .out(SD48));
lcell U48(.in(SD48)  , .out(SD49));
lcell U49(.in(SD49)  , .out(SD50));
lcell U50(.in(SD50)  , .out(SD51));
lcell U51(.in(SD51)  , .out(SD52));
lcell U52(.in(SD52)  , .out(SD53));
lcell U53(.in(SD53)  , .out(SD54));
lcell U54(.in(SD54)  , .out(SD55));
lcell U55(.in(SD55)  , .out(SD56));
lcell U56(.in(SD56)  , .out(SD57));
lcell U57(.in(SD57)  , .out(SD58));
lcell U58(.in(SD58)  , .out(SD59));
lcell U59(.in(SD59)  , .out(SD60));
lcell U60(.in(SD60)  , .out(SD61));
lcell U61(.in(SD61)  , .out(SD62));
lcell U62(.in(SD62)  , .out(SD63));
lcell U63(.in(SD63)  , .out(SD64));
lcell U64(.in(SD64)  , .out(SD65));
lcell U65(.in(SD65)  , .out(SD66));
lcell U66(.in(SD66)  , .out(SD67));
lcell U67(.in(SD67)  , .out(SD68));
lcell U68(.in(SD68)  , .out(SD69));
lcell U69(.in(SD69)  , .out(SD70));
lcell U70(.in(SD70)  , .out(SD71));
lcell U71(.in(SD71)  , .out(SD72));
lcell U72(.in(SD72)  , .out(SD73));
lcell U73(.in(SD73)  , .out(SD74));
lcell U74(.in(SD74)  , .out(SD75));
lcell U75(.in(SD75)  , .out(SD76));
lcell U76(.in(SD76)  , .out(SD77));
lcell U77(.in(SD77)  , .out(SD78));
lcell U78(.in(SD78)  , .out(SD79));
lcell U79(.in(SD79)  , .out(D80));

endmodule
