module DLY_chain(
    IN,
    D80,
);

input   IN;
output  D80;

lcell  U0/* synthesis keep */(.in(IN)    , .out(SD1));
lcell  U1/* synthesis keep */(.in(SD1)   , .out(SD2));
lcell  U2/* synthesis keep */(.in(SD2)   , .out(SD3));
lcell  U3/* synthesis keep */(.in(SD3)   , .out(SD4));
lcell  U4/* synthesis keep */(.in(SD4)   , .out(SD5));
lcell  U5/* synthesis keep */(.in(SD5)   , .out(SD6));
lcell  U6/* synthesis keep */(.in(SD6)   , .out(SD7));
lcell  U7/* synthesis keep */(.in(SD7)   , .out(SD8));
lcell  U8/* synthesis keep */(.in(SD8)   , .out(SD9));
lcell  U9/* synthesis keep */(.in(SD9)   , .out(SD10));
lcell U10/* synthesis keep */(.in(SD10)  , .out(SD11));
lcell U11/* synthesis keep */(.in(SD11)  , .out(SD12));
lcell U12/* synthesis keep */(.in(SD12)  , .out(SD13));
lcell U13/* synthesis keep */(.in(SD13)  , .out(SD14));
lcell U14/* synthesis keep */(.in(SD14)  , .out(SD15));
lcell U15/* synthesis keep */(.in(SD15)  , .out(SD16));
lcell U16/* synthesis keep */(.in(SD16)  , .out(SD17));
lcell U17/* synthesis keep */(.in(SD17)  , .out(SD18));
lcell U18/* synthesis keep */(.in(SD18)  , .out(SD19));
lcell U19/* synthesis keep */(.in(SD19)  , .out(SD20));
lcell U20/* synthesis keep */(.in(SD20)  , .out(SD21));
lcell U21/* synthesis keep */(.in(SD21)  , .out(SD22));
lcell U22/* synthesis keep */(.in(SD22)  , .out(SD23));
lcell U23/* synthesis keep */(.in(SD23)  , .out(SD24));
lcell U24/* synthesis keep */(.in(SD24)  , .out(SD25));
lcell U25/* synthesis keep */(.in(SD25)  , .out(SD26));
lcell U26/* synthesis keep */(.in(SD26)  , .out(SD27));
lcell U27/* synthesis keep */(.in(SD27)  , .out(SD28));
lcell U28/* synthesis keep */(.in(SD28)  , .out(SD29));
lcell U29/* synthesis keep */(.in(SD29)  , .out(SD30));
lcell U30/* synthesis keep */(.in(SD30)  , .out(SD31));
lcell U31/* synthesis keep */(.in(SD31)  , .out(SD32));
lcell U32/* synthesis keep */(.in(SD32)  , .out(SD33));
lcell U33/* synthesis keep */(.in(SD33)  , .out(SD34));
lcell U34/* synthesis keep */(.in(SD34)  , .out(SD35));
lcell U35/* synthesis keep */(.in(SD35)  , .out(SD36));
lcell U36/* synthesis keep */(.in(SD36)  , .out(SD37));
lcell U37/* synthesis keep */(.in(SD37)  , .out(SD38));
lcell U38/* synthesis keep */(.in(SD38)  , .out(SD39));
lcell U39/* synthesis keep */(.in(SD39)  , .out(SD40));
lcell U40/* synthesis keep */(.in(SD40)  , .out(SD41));
lcell U41/* synthesis keep */(.in(SD41)  , .out(SD42));
lcell U42/* synthesis keep */(.in(SD42)  , .out(SD43));
lcell U43/* synthesis keep */(.in(SD43)  , .out(SD44));
lcell U44/* synthesis keep */(.in(SD44)  , .out(SD45));
lcell U45/* synthesis keep */(.in(SD45)  , .out(SD46));
lcell U46/* synthesis keep */(.in(SD46)  , .out(SD47));
lcell U47/* synthesis keep */(.in(SD47)  , .out(SD48));
lcell U48/* synthesis keep */(.in(SD48)  , .out(SD49));
lcell U49/* synthesis keep */(.in(SD49)  , .out(SD50));
lcell U50/* synthesis keep */(.in(SD50)  , .out(SD51));
lcell U51/* synthesis keep */(.in(SD51)  , .out(SD52));
lcell U52/* synthesis keep */(.in(SD52)  , .out(SD53));
lcell U53/* synthesis keep */(.in(SD53)  , .out(SD54));
lcell U54/* synthesis keep */(.in(SD54)  , .out(SD55));
lcell U55/* synthesis keep */(.in(SD55)  , .out(SD56));
lcell U56/* synthesis keep */(.in(SD56)  , .out(SD57));
lcell U57/* synthesis keep */(.in(SD57)  , .out(SD58));
lcell U58/* synthesis keep */(.in(SD58)  , .out(SD59));
lcell U59/* synthesis keep */(.in(SD59)  , .out(SD60));
lcell U60/* synthesis keep */(.in(SD60)  , .out(SD61));
lcell U61/* synthesis keep */(.in(SD61)  , .out(SD62));
lcell U62/* synthesis keep */(.in(SD62)  , .out(SD63));
lcell U63/* synthesis keep */(.in(SD63)  , .out(SD64));
lcell U64/* synthesis keep */(.in(SD64)  , .out(SD65));
lcell U65/* synthesis keep */(.in(SD65)  , .out(SD66));
lcell U66/* synthesis keep */(.in(SD66)  , .out(SD67));
lcell U67/* synthesis keep */(.in(SD67)  , .out(SD68));
lcell U68/* synthesis keep */(.in(SD68)  , .out(SD69));
lcell U69/* synthesis keep */(.in(SD69)  , .out(SD70));
lcell U70/* synthesis keep */(.in(SD70)  , .out(SD71));
lcell U71/* synthesis keep */(.in(SD71)  , .out(SD72));
lcell U72/* synthesis keep */(.in(SD72)  , .out(SD73));
lcell U73/* synthesis keep */(.in(SD73)  , .out(SD74));
lcell U74/* synthesis keep */(.in(SD74)  , .out(SD75));
lcell U75/* synthesis keep */(.in(SD75)  , .out(SD76));
lcell U76/* synthesis keep */(.in(SD76)  , .out(SD77));
lcell U77/* synthesis keep */(.in(SD77)  , .out(SD78));
lcell U78/* synthesis keep */(.in(SD78)  , .out(SD79));
lcell U79/* synthesis keep */(.in(SD79)  , .out(D80));

endmodule
